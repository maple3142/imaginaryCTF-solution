module sat(out, in);
    input [255:0] in;
    output out;

or(o88, in[235], ~in[236], ~in[237]);
and(o79, in[211], in[212], in[213]);
or(o85, in[227], in[228], ~in[229]);
and(t13, t6, t7, t8);
and(t7, r21, r22, r23);
or(o51, ~in[136], in[137], in[138]);
and(o84, ~in[224], in[225], in[226]);
and(o4, ~in[11], in[12], in[13]);
and(t9, r27, r28, r29);
and(t11, t0, t1, t2);
and(t1, r3, r4, r5);
and(r28, o84, ~o85, o86);
and(o31, in[83], ~in[84], in[85]);
and(o1, in[3], in[4], in[5]);
and(r21, ~o63, o64, ~o65);
or(o69, ~in[184], ~in[185], ~in[186]);
and(o42, in[112], in[113], in[114]);
or(o44, ~in[118], in[119], ~in[118]);
or(o57, ~in[152], in[153], in[154]);
and(r31, o93, ~o94, ~o95);
and(r3, ~o9, ~o10, ~o11);
and(o29, in[78], ~in[79], in[78]);
and(t8, r24, r25, r26);
and(o64, ~in[171], in[172], in[173]);
or(o23, ~in[62], in[63], ~in[62]);
or(o55, in[147], in[148], ~in[149]);
or(o60, in[160], in[161], ~in[162]);
and(o93, in[248], ~in[249], ~in[250]);
and(r15, ~o45, o46, o47);
or(o59, ~in[158], in[159], ~in[158]);
and(r4, o12, o13, o14);
or(o90, ~in[240], ~in[241], in[242]);
and(r18, ~o54, ~o55, o56);
and(o62, in[166], ~in[167], in[166]);
or(o45, in[120], in[121], ~in[122]);
and(o35, in[94], ~in[95], in[94]);
or(o80, in[214], in[215], in[214]);
and(o30, ~in[80], in[81], in[82]);
and(r29, o87, ~o88, o89);
and(o41, in[110], ~in[111], in[110]);
and(o49, ~in[131], in[132], in[133]);
and(t6, r18, r19, r20);
or(o63, in[168], in[169], in[170]);
or(o81, ~in[216], ~in[217], in[218]);
and(o89, in[238], ~in[239], in[238]);
or(o18, ~in[48], ~in[49], ~in[50]);
or(o37, ~in[99], in[100], ~in[101]);
and(t12, t3, t4, t5);
and(o38, in[102], ~in[103], in[102]);
and(r23, ~o69, o70, o71);
and(o71, in[190], ~in[191], in[190]);
and(o14, in[38], ~in[39], in[38]);
or(o58, ~in[155], in[156], ~in[157]);
and(r19, ~o57, ~o58, ~o59);
and(o47, in[126], ~in[127], in[126]);
or(o52, in[139], in[140], ~in[141]);
and(r27, ~o81, ~o82, ~o83);
or(o28, ~in[75], ~in[76], in[77]);
and(o17, in[46], ~in[47], in[46]);
or(o61, ~in[163], in[164], ~in[165]);
and(r7, o21, o22, ~o23);
or(o40, in[107], ~in[108], ~in[109]);
or(o16, in[43], ~in[44], ~in[45]);
and(r13, ~o39, ~o40, o41);
and(o86, in[230], ~in[231], in[230]);
or(o50, ~in[134], in[135], ~in[134]);
and(o46, ~in[123], ~in[124], in[125]);
and(o8, in[22], ~in[23], in[22]);
or(o33, ~in[88], in[89], in[90]);
or(o66, ~in[176], in[177], ~in[178]);
or(o73, in[195], in[196], ~in[197]);
and(t5, r15, r16, r17);
and(o12, in[32], ~in[33], in[34]);
and(o87, ~in[232], ~in[233], in[234]);
or(o67, ~in[179], in[180], ~in[181]);
and(r0, o0, o1, o2);
and(t3, r9, r10, r11);
and(t10, r30, r31, r17);
or(o92, ~in[246], in[247], ~in[246]);
and(t2, r6, r7, r8);
or(o54, ~in[144], ~in[145], in[146]);
and(o72, in[192], in[193], ~in[194]);
and(r2, ~o6, ~o7, o8);
and(o0, in[0], ~in[1], in[2]);
and(r5, o15, ~o16, o17);
or(o94, ~in[251], in[252], ~in[253]);
and(r30, ~o90, o91, ~o92);
and(r17, ~o51, ~o52, o53);
and(out, t12, t13, t14);
and(r6, ~o18, o19, ~o20);
and(o56, in[150], ~in[151], in[150]);
and(r11, ~o33, ~o34, o35);
and(o53, in[142], ~in[143], in[142]);
and(r9, ~o27, ~o28, o29);
or(o27, ~in[72], ~in[73], ~in[74]);
and(o24, in[64], ~in[65], ~in[66]);
and(t0, r0, r1, r2);
or(o6, ~in[16], in[17], ~in[18]);
and(o68, in[182], ~in[183], in[182]);
and(r24, o72, ~o73, o74);
and(o74, in[198], ~in[199], in[198]);
and(r10, o30, o31, ~o32);
and(o25, in[67], ~in[68], in[69]);
or(o11, ~in[30], in[31], ~in[30]);
or(o32, ~in[86], in[87], ~in[86]);
or(o82, ~in[219], ~in[220], ~in[221]);
or(o9, ~in[24], in[25], ~in[26]);
and(o43, in[115], in[116], ~in[117]);
and(o78, ~in[208], ~in[209], in[210]);
or(o77, ~in[206], in[207], ~in[206]);
and(o19, in[51], in[52], ~in[53]);
or(o20, ~in[54], in[55], ~in[54]);
or(o7, ~in[19], in[20], ~in[21]);
and(t14, t9, t10, t11);
and(o13, ~in[35], ~in[36], in[37]);
and(o21, ~in[56], ~in[57], in[58]);
and(r16, ~o48, o49, ~o50);
and(o22, ~in[59], in[60], in[61]);
and(o5, in[14], ~in[15], in[14]);
and(o91, ~in[243], ~in[244], in[245]);
and(r26, o78, o79, ~o80);
or(o83, ~in[222], in[223], ~in[222]);
or(o3, ~in[8], ~in[9], in[10]);
or(o75, ~in[200], ~in[201], ~in[202]);
and(r14, o42, o43, ~o44);
or(o95, ~in[254], in[255], ~in[254]);
or(o34, in[91], in[92], ~in[93]);
and(r25, ~o75, o76, ~o77);
and(o26, in[70], ~in[71], in[70]);
and(t4, r12, r13, r14);
and(r22, ~o66, ~o67, o68);
and(r12, ~o36, ~o37, o38);
and(o2, in[6], ~in[7], in[6]);
or(o39, in[104], in[105], ~in[106]);
and(r20, ~o60, ~o61, o62);
or(o36, in[96], in[97], in[98]);
and(r8, o24, o25, o26);
and(o76, in[203], in[204], ~in[205]);
or(o65, ~in[174], in[175], ~in[174]);
or(o10, in[27], in[28], ~in[29]);
and(o70, in[187], ~in[188], in[189]);
and(r1, ~o3, o4, o5);
or(o48, in[128], in[129], ~in[130]);
and(o15, in[40], in[41], ~in[42]);

endmodule

module main;
    wire [255:0] flag = 256'h696374667b00000000000000000000000000000000000000000000000000007d;
    wire valid;

    sat flagchecker(valid, flag);

    initial begin
        #50;
        if (valid) begin
            $display("Correct!");
            $finish;
        end
        $display("Incorrect flag...");
    end
endmodule